../II_full/ntt_addr_gen.vhd