../II_sign/double_bfu.vhd