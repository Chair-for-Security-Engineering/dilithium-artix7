../II_verify/keccak_round.vhd