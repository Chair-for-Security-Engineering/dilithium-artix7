../II_sign/macc_poly.vhd