../II_sign/keccak.vhd