../II_verify/red_dsp_3.vhd