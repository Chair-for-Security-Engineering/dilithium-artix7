../II_verify/sign.vhd