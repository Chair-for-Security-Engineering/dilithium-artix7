../II_verify/ntt_addr_gen.vhd