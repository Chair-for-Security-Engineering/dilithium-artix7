../II_full/reg32.vhd