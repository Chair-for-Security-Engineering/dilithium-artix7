../II_full/dyn_shift_reg.vhd