../II_verify/bfu_adder.vhd