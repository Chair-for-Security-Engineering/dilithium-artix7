../II_full/use_hint_lut.vhd