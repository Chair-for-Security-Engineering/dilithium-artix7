../II_verify/expand_y.vhd