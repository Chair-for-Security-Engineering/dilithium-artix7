../II_verify/mem_8_poly.vhd