../II_verify/bfu_reducer.vhd