../II_full/hreg.vhd