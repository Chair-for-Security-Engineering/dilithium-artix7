../II_sign/red_dsp.vhd