../II_full/parmset.vhd