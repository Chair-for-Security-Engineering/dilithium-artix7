../II_sign/butterfly_dsp.vhd