../II_full/macc_coeff.vhd