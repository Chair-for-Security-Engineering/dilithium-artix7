../II_sign/convert_yz.vhd