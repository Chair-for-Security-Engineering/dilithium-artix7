../II_verify/reg32.vhd