../II_verify/macc_coeff.vhd