../II_sign/memory.vhd