../II_full/sample_y_dsp.vhd