../II_sign/keccak_counter.vhd