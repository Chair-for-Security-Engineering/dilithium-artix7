../II_sign/red_dsp_2.vhd