../II_sign/store.vhd