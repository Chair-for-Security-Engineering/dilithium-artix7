../II_verify/keccak_settings.vhd