../II_sign/hreg.vhd