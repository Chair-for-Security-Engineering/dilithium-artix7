../II_full/red_dsp_1.vhd