../II_verify/keccak_controller.vhd