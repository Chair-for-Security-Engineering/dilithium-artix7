../II_verify/keccak_rc.vhd