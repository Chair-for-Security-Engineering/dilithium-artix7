../II_verify/digest_msg.vhd