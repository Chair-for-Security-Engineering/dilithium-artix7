../II_sign/mem_8_poly.vhd