../II_sign/expand_y.vhd