../II_sign/ntt.vhd