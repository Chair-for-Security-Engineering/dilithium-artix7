../II_sign/use_hint.vhd