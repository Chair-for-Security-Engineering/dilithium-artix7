../II_verify/macc_poly.vhd