../II_sign/unpack_yz.vhd