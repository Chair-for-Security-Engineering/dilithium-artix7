../II_full/ntt.vhd