../II_sign/keccak_settings.vhd