../II_verify/counter.vhd