../II_full/keccak_settings.vhd