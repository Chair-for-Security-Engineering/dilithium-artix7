../II_full/mem_8_poly.vhd