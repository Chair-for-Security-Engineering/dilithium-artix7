../II_verify/globals.vhd