../II_full/verify.vhd