../II_verify/keygen.vhd