../II_sign/red_dsp_1.vhd