../II_verify/bfu_subtractor.vhd