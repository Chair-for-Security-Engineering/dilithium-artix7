../II_full/unpack_yz.vhd