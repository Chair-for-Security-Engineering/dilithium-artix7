../II_verify/red_dsp_2.vhd