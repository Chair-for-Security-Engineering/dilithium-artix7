../II_verify/interfaces.vhd