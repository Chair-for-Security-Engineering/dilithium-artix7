../II_sign/sign.vhd