../II_sign/verify_precomp.vhd