../II_sign/load.vhd