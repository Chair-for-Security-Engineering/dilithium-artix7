../II_sign/bfu_adder.vhd