../II_verify/check_z.vhd