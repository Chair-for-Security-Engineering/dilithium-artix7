../II_verify/hreg.vhd