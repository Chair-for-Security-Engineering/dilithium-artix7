../II_verify/sign_precomp.vhd