../II_verify/use_hint.vhd