../II_verify/keccak.vhd