../II_full/bfu_adder.vhd