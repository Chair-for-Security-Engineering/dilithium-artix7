../II_verify/bfu_stage_2.vhd