../II_sign/ntt_addr_gen.vhd