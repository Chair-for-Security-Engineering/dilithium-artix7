../II_full/expand.vhd