../II_full/keccak_rc.vhd