../II_full/sign.vhd