../II_sign/ballsample.vhd