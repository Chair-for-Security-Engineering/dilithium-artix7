../II_verify/crh_rho_t1.vhd