../II_full/red_dsp.vhd