../II_sign/highbits.vhd