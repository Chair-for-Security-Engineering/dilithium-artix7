../V_full/parmset.vhd