../II_sign/bfu_subtractor.vhd