../II_full/interfaces.vhd