../II_full/sign_precomp.vhd