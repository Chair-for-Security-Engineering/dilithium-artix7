../II_full/double_bfu.vhd