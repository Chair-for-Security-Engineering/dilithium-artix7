../II_verify/butterfly_dsp.vhd