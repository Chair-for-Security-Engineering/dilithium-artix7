../II_sign/check_z.vhd