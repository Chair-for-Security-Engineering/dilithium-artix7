../II_sign/macc_coeff.vhd