../II_verify/expand.vhd