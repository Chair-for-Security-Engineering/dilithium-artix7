../II_full/keccak_controller.vhd