../II_full/bfu_stage_1.vhd