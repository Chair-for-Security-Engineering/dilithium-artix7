../II_verify/convert_yz.vhd