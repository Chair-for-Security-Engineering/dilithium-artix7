../II_verify/load.vhd