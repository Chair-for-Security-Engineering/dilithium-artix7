../II_full/bfu_stage_2.vhd