../II_sign/reg32.vhd