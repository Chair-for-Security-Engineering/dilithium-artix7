../II_sign/digest_msg.vhd