../II_sign/mem_8_quarter_poly.vhd