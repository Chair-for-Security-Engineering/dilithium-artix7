../II_sign/keccak_round.vhd