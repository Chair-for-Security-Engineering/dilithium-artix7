../II_full/check_z.vhd