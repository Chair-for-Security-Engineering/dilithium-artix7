../II_sign/keygen.vhd