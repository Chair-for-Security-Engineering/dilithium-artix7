../II_verify/store.vhd