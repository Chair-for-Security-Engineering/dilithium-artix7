../II_sign/globals.vhd