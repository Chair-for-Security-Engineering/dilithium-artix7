../II_sign/macc_dsp.vhd