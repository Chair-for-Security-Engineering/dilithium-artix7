../II_sign/red_dsp_3.vhd