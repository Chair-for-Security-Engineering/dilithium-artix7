../II_full/keccak.vhd