../II_verify/ballsample.vhd