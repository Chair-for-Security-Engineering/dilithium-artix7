../II_full/expands1s2.vhd