../II_verify/red_dsp.vhd