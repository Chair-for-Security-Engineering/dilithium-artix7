../II_sign/use_hint_lut.vhd