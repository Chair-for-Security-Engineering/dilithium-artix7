../II_verify/dyn_shift_reg.vhd