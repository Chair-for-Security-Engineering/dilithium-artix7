../II_verify/expands1s2.vhd