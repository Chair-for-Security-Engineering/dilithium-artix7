../II_sign/keccak_controller.vhd