../II_full/counter.vhd