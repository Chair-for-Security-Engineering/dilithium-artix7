../II_verify/use_hint_lut.vhd