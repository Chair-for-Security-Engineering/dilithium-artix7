../II_verify/ntt.vhd