../II_sign/matmul.vhd