../II_full/convert_yz.vhd