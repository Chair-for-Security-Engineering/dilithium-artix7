../II_full/globals.vhd