../II_sign/bfu_reducer.vhd