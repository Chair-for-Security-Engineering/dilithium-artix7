../II_verify/keccak_counter.vhd