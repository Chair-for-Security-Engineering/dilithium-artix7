../II_verify/verify.vhd