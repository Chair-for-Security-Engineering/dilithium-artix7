../II_sign/sign_precomp.vhd