../II_full/digest_msg.vhd