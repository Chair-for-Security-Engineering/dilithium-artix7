../II_full/use_hint.vhd