../II_full/store.vhd