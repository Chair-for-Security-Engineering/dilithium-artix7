../II_sign/expands1s2.vhd