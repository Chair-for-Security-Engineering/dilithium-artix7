../II_full/red_dsp_2.vhd