../II_sign/keccak_rc.vhd