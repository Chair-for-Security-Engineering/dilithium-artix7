../II_sign/counter.vhd