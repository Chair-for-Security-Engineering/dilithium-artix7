../II_full/macc_poly.vhd