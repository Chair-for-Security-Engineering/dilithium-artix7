../II_verify/red_dsp_1.vhd