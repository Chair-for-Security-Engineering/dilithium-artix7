../II_full/load.vhd