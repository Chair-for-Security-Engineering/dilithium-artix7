../II_full/memory.vhd