../II_verify/memory.vhd