../II_sign/bfu_stage_1.vhd