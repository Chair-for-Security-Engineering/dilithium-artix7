../II_full/ballsample.vhd