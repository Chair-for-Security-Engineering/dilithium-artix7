../II_sign/sample_y_dsp.vhd