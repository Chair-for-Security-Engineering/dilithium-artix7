../II_full/keccak_counter.vhd