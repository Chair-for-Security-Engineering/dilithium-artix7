../II_verify/double_bfu.vhd