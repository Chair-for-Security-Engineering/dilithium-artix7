../II_sign/bfu_stage_2.vhd