../II_full/crh_rho_t1.vhd