../II_full/verify_precomp.vhd