../II_sign/verify.vhd