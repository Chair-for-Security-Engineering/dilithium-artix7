../II_verify/sample_y_dsp.vhd