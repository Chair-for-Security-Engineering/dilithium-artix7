../II_verify/matmul.vhd