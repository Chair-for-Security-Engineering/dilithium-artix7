../II_sign/dilithium_top.vhd