../II_sign/crh_rho_t1.vhd