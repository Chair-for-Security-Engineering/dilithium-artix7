../II_full/mem_8_quarter_poly.vhd