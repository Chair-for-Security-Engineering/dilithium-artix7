../II_sign/red_dsp_4.vhd