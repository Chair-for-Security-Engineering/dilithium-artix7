../II_sign/mem_twiddle.vhd