../II_full/mem_twiddle.vhd