../II_verify/highbits2gamma.vhd