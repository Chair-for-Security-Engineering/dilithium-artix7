../II_full/expand_y.vhd