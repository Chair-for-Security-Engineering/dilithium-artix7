../II_verify/mem_8_quarter_poly.vhd