../II_verify/dilithium_top.vhd