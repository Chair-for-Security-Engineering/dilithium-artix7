../II_full/keygen.vhd