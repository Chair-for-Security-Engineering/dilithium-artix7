../II_sign/interfaces.vhd