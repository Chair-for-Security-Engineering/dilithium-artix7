../II_verify/highbits.vhd