../II_full/dilithium_top.vhd