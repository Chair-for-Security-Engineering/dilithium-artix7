../II_full/keccak_round.vhd