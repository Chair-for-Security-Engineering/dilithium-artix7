../II_verify/macc_dsp.vhd