../II_verify/verify_precomp.vhd