../II_verify/mem_twiddle.vhd