../II_sign/dyn_shift_reg.vhd