../II_sign/expand.vhd