../II_sign/highbits2gamma.vhd