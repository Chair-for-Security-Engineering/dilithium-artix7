../II_verify/unpack_yz.vhd