../II_verify/red_dsp_4.vhd