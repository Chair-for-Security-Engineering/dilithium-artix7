../II_verify/bfu_stage_1.vhd